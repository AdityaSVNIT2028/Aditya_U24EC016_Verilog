`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: SVNIT
// Engineer: Aditya
//////////////////////////////////////////////////////////////////////////////////

module mux_2X1(input i0, i1, i_s,
output reg Y
    );
    always @(*) begin
    if(!i_s)
    Y = i0;
    else
    Y = i1;
    end
endmodule
